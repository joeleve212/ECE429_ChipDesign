*** SPICE deck for cell test_inv1{sch} from library White_inverters
*** Created on Tue Feb 04, 2014 11:19:28
*** Last revised on Sun Feb 02, 2020 23:52:52
*** Written on Mon Feb 10, 2020 09:56:18 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT White_inverters__inv1 FROM CELL inv1{sch}
.SUBCKT White_inverters__inv1 in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd N L=0.6U W=1.2U
Mpmos@0 vdd in out vdd P L=0.6U W=1.2U
.ENDS White_inverters__inv1

.global gnd vdd

*** TOP LEVEL CELL: test_inv1{sch}
VPulse@1 a0 gnd DC=0 pulse 0 5 0ns 10p 10p 0.5n 1n
Xinv1@0 a0 a1 White_inverters__inv1
Xinv1@1 a1 a2 White_inverters__inv1
Xinv1@2 a2 a3 White_inverters__inv1

* Spice Code nodes in cell cell 'test_inv1{sch}'
.tran 2n
.meas tran tpHL trig v(a1) val=2.5 rise=1 targ v(a2) val=2.5 fall=1
.meas tran tpLH trig v(a1) val=2.5 fall=1 targ v(a2) val=2.5 rise=1
.meas tran tpavg param (tpHL+tpLH)/2
.meas tran trise trig v(a2) val='0.10*5' rise=1 targ v(a2) val='0.90*5' rise=1
.meas tran tfall trig v(a2) val='0.90*5' fall=1 targ v(a2) val='0.10*5' fall=1
Vdd vdd 0 5
Vgd gnd 0 0
.include c5.txt
.END
