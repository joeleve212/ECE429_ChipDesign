*** SPICE deck for cell test_Cell{sch} from library Leveille_HW7
*** 
*** ECE 429
*** Valparaiso University
*** 
*** Project settings version ** 3 **
*** 
*** Created on Wed Mar 25, 2020 17:41:12
*** Last revised on Wed Mar 25, 2020 18:13:34
*** Written on Wed Mar 25, 2020 18:14:29 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Leveille_HW7__inv FROM CELL Leveille_HW7:inv{sch}
.SUBCKT Leveille_HW7__inv x y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 y x gnd gnd N L=0.6U W=1.8U
Mpmos@0 vdd x y vdd P L=0.6U W=3U
.ENDS Leveille_HW7__inv

*** SUBCIRCUIT Leveille_HW7__transGate FROM CELL Leveille_HW7:transGate{sch}
.SUBCKT Leveille_HW7__transGate CLK in inv_CLK out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out CLK in gnd N L=0.6U W=0.6U
Mpmos@0 in inv_CLK out vdd P L=0.6U W=0.6U
.ENDS Leveille_HW7__transGate

*** SUBCIRCUIT Leveille_HW7__D_latch FROM CELL Leveille_HW7:D_latch{sch}
.SUBCKT Leveille_HW7__D_latch clk D D_out inv_clk inv_D
** GLOBAL gnd
** GLOBAL vdd
Xinv@2 D_out inv_D Leveille_HW7__inv
Xinv@3 inv_D net@41 Leveille_HW7__inv
XtransGat@1 clk D inv_clk D_out Leveille_HW7__transGate
XtransGat@2 inv_clk net@41 clk D_out Leveille_HW7__transGate
.ENDS Leveille_HW7__D_latch

*** SUBCIRCUIT Leveille_HW7__D_FF FROM CELL Leveille_HW7:D_FF{sch}
.SUBCKT Leveille_HW7__D_FF /clk /Q clk D Q
** GLOBAL gnd
** GLOBAL vdd
XD_latch@0 /clk net@0 D_latch@0_D_out clk net@2 Leveille_HW7__D_latch
XD_latch@1 clk net@2 net@27 /clk net@5 Leveille_HW7__D_latch
Xinv@0 D net@0 Leveille_HW7__inv
Xinv@1 net@27 /Q Leveille_HW7__inv
Xinv@2 net@5 Q Leveille_HW7__inv
.ENDS Leveille_HW7__D_FF

.global gnd vdd

*** TOP LEVEL CELL: Leveille_HW7:test_Cell{sch}
XD_FF@0 ckb Qbar ck rd Q Leveille_HW7__D_FF
Xinv@0 D net@9 Leveille_HW7__inv
Xinv@1 CLK ckb Leveille_HW7__inv
Xinv@2 ckb ck Leveille_HW7__inv
Xinv@4 net@9 rd Leveille_HW7__inv
Xinv@8 Qbar OUT Leveille_HW7__inv
Xinv@9 Qbar OUT Leveille_HW7__inv
Xinv@10 Qbar OUT Leveille_HW7__inv
Xinv@11 Qbar OUT Leveille_HW7__inv
Xinv@12 Q OUT Leveille_HW7__inv
Xinv@13 Q OUT Leveille_HW7__inv
Xinv@14 Q OUT Leveille_HW7__inv
Xinv@15 Q OUT Leveille_HW7__inv

* Spice Code nodes in cell cell 'Leveille_HW7:test_Cell{sch}'
VGND GND 0 DC 0
VVDD VDD 0 DC 5
VCLK CLK 0 DC 0 PULSE 0 5 0 10p 10p 3n 6n
VIN D 0 DC 0 PULSE 5 0 200p 10p 10p 3n 5.99n
.include c5.txt
.tran 2000n UIC
.save v(rd) v(ck) v(q) v(qbar) v(D_FF@2:D_latch@0:x) v(D_FF@2:outbar) v(D_FF@2:D_latch@1:x) v(D_FF@2:mid) dialogbox
*.options post
.END
