*** SPICE deck for cell inv2{sch} from library Leveille_hw5
*** Created on Wed Feb 19, 2020 11:48:42
*** Last revised on Wed Feb 19, 2020 12:06:48
*** Written on Thu Feb 20, 2020 15:16:36 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: inv2{sch}
Mnmos@0 y Vin gnd gnd NMOS L=0.6U W=7.2U
Mpmos@0 vdd Vin y vdd PMOS L=0.6U W=14.4U

* Spice Code nodes in cell cell 'inv2{sch}'
Vdd vdd 0 5
Vgd gnd 0 0
.include c5.txt
.END
